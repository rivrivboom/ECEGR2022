--------------------------------------------------------------------------------
--
-- Test Bench for LAB #4
--
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;

ENTITY testALU_vhd IS
END testALU_vhd;

ARCHITECTURE behavior OF testALU_vhd IS 

	-- Component Declaration for the Unit Under Test (UUT)
	COMPONENT ALU
		Port(	DataIn1: in std_logic_vector(31 downto 0);
			DataIn2: in std_logic_vector(31 downto 0);
			ALUCtrl: in std_logic_vector(4 downto 0);
			Zero: out std_logic;
			ALUResult: out std_logic_vector(31 downto 0) );
	end COMPONENT ALU;

	--Inputs
	SIGNAL datain_a : std_logic_vector(31 downto 0) := (others=>'0');
	SIGNAL datain_b : std_logic_vector(31 downto 0) := (others=>'0');
	SIGNAL control	: std_logic_vector(4 downto 0)	:= (others=>'0');

	--Outputs
	SIGNAL result   :  std_logic_vector(31 downto 0);
	SIGNAL zeroOut  :  std_logic;

BEGIN

	-- Instantiate the Unit Under Test (UUT)
	uut: ALU PORT MAP(
		DataIn1 => datain_a,
		DataIn2 => datain_b,
		ALUCtrl => control,
		Zero => zeroOut,
		ALUResult => result
	);
	

	tb : PROCESS
BEGIN

		-- Wait 100 ns for global reset to finish
		wait for 100 ns;

		-- Start testing the ALU

		--add
		control  <= "0000X";	
		datain_a <= X"01234567";	-- DataIn in hex
		datain_b <= X"11223344";

		--result;	-- Control in binary )
		
		wait for 20 ns; 			

		--sub
		datain_a <= X"ABABABAB";	-- DataIn in hex
		datain_b <= X"11223344";
		control  <= "0001X";		-- Control in binary
		
		wait for 20 ns; 			

	 			
		--and
		datain_b <= X"FFFFFFFF" ;	-- DataIn in binary
		control  <= "0010X";		-- Control in binary 
		
		wait for 20 ns; 			

		

		--or
		datain_a <= X"11110011";	-- DataIn in binary
		datain_b <= X"11001100";
		control  <= "011XX";		-- Control in binary 
		
		wait for 20 ns; 			


		--sll
		datain_a <= X"CBACBDFF";	-- DataIn in hex
		datain_b <= X"00000002";
		control  <= "0010X";		-- Control in binary
		
		wait for 20 ns; 			-- result = 0x00000008  and zeroOut = 0


		--srl
		control  <= "0011X";		-- Control in binary 
		
		wait for 20 ns; 			-- result = 0x00000001  and zeroOut = 0

		control <= "1XXXX";
		wait for 20 ns; 			-- result = 0x00000001  and zeroOut = 0

		wait;
	end process;
end;
